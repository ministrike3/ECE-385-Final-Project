// The point of this code is to decide whether or not to print the protagonist
// Neil, in his regular or powered form.

// he becomes powered when he eats the 4th coin that appears on the screen
// which represents the change from TTL to Verilog!

// The module works by taking a signal called power that changes from 0 to 1
// when the hero sprite onscreen collides with the powerup coin
// that changes the internal signal called change from 0 to 1 in this module.

// the middle of the code declares 2 sprite arrays, powerhero and hero123.

// At the bottom, an always comb loop decides (based on if change = 1 or 0)
// to declare the output hero_text
// to equal either powerhero or hero123.


module hero_sprite_decider(
									input logic clk,
									input power,
									output logic [0:79][0:39][0:5] hero_text
									);

logic [0:79][0:39][0:5] powerhero_text;
logic [0:79][0:39][0:5] hero123_text;

logic change = 0;
always_ff@(posedge clk)
begin
	if ((change==0)&&(power==1))
	begin
	change<=1;
	end
	else
	change<=change;

end


always_comb
begin
hero123_text <=
//hero_text <=
'{
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,42,2,1,45,46,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,42,2,1,45,46,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,1,46,43,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,46,46,46,45,1,1,1,42,15,46,46,46,46,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,46,45,46,46,46,42,45,1,1,1,42,15,46,45,46,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,43,46,2,2,15,42,1,1,1,2,2,42,43,46,46,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,2,1,15,42,1,2,15,43,46,2,1,1,1,43,43,46,46,46,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,2,2,15,42,1,1,46,46,46,2,1,1,1,43,43,46,46,46,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,46,42,15,46,1,1,1,2,2,46,2,1,1,45,46,43,46,45,2,2,43,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,46,42,15,46,1,1,1,1,2,42,2,1,1,1,46,15,42,46,1,1,15,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,45,46,15,46,1,1,1,1,2,46,2,1,1,1,46,15,42,46,1,2,43,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,1,2,15,43,42,45,43,43,43,15,42,1,2,15,42,1,2,15,43,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,1,2,15,15,42,46,15,15,15,15,42,1,2,24,43,1,2,15,15,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,2,2,43,43,42,46,43,43,43,43,43,2,2,2,45,1,45,15,43,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,43,43,15,43,45,42,15,23,21,36,36,36,36,21,23,1,2,46,43,15,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,15,15,15,43,13,42,15,23,21,36,36,36,36,21,23,1,2,13,43,15,42,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,43,43,43,43,23,23,43,36,21,36,22,22,36,21,36,43,23,23,43,43,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,45,42,46,23,21,21,21,36,36,20,7,7,20,36,21,21,21,21,23,45,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,45,42,13,46,21,36,36,36,36,20,7,7,20,36,36,36,36,21,46,13,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,43,46,46,23,23,21,36,36,36,12,4,4,4,12,12,36,36,36,21,23,23,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,46,46,21,21,36,36,36,12,20,37,15,45,43,20,12,36,36,36,21,21,46,45,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,43,46,46,36,36,36,21,21,12,20,37,19,45,43,20,12,21,21,36,36,36,46,13,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,43,2,2,36,36,21,36,19,35,12,12,12,12,12,12,35,19,36,21,36,36,2,2,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,46,46,45,43,43,1,1,36,36,21,19,35,35,35,4,20,20,4,35,35,35,19,21,36,36,1,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,46,46,45,42,42,1,1,21,21,21,24,35,35,35,4,20,20,4,35,35,35,19,21,21,21,1,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,33,39,45,2,2,2,35,35,35,35,35,35,35,35,35,35,35,35,35,35,2,2,2,45,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,40,38,42,45,1,2,35,35,35,35,35,35,35,35,35,35,35,35,35,35,2,1,45,42,41,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,33,40,42,45,1,2,35,35,35,35,35,35,35,35,35,35,35,35,35,35,2,1,45,42,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,39,39,45,45,33,41,3,12,2,42,42,42,42,42,42,42,42,2,12,3,41,33,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,40,45,45,39,38,7,12,1,2,45,45,45,45,45,45,2,1,12,7,38,39,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,39,45,45,39,38,7,12,1,45,45,45,45,45,45,45,45,1,12,7,48,39,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,55,55,7,12,1,37,55,54,54,54,54,55,37,1,12,3,55,55,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,55,5,7,12,1,37,55,54,55,55,54,55,37,1,12,7,55,55,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,54,55,3,12,2,47,55,54,54,54,54,55,37,2,12,3,54,54,2,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,45,45,1,43,55,54,55,55,55,55,54,54,54,55,54,54,54,54,42,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,45,45,2,15,55,55,55,55,54,55,55,55,55,54,54,54,54,55,15,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,42,38,38,38,54,55,38,38,38,38,55,54,38,48,38,42,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,1,1,45,44,48,55,33,44,44,33,55,48,44,45,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,1,1,42,39,38,55,39,44,44,39,55,38,39,42,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,42,42,23,23,15,24,37,15,15,15,15,37,24,15,23,23,42,42,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,2,35,35,22,36,1,1,1,2,45,45,2,1,1,1,36,22,35,35,46,2,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,35,35,22,36,1,1,1,45,46,13,45,1,1,1,36,22,35,35,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,24,37,19,43,23,23,19,23,21,19,19,36,36,43,43,36,23,23,36,12,37,33,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,1,1,38,38,23,23,1,42,35,36,22,35,35,22,22,35,35,22,23,1,21,22,54,38,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,1,1,1,40,38,23,23,1,43,35,36,22,35,35,22,22,35,35,22,23,1,21,22,54,38,1,1,1,0,0,0,0,0,0},
'{0,0,0,0,0,24,54,33,15,47,48,2,2,0,0,42,19,35,36,36,35,35,22,36,23,0,0,23,23,38,38,33,33,54,24,0,0,0,0,0},
'{0,0,0,0,1,37,6,48,39,47,48,2,0,0,0,1,19,35,22,22,35,35,22,21,1,0,0,0,2,38,38,48,38,6,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,40,39,48,48,2,0,0,0,1,19,35,22,22,35,35,22,21,1,0,0,0,2,38,38,39,47,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,55,55,42,2,0,0,2,2,1,36,22,35,35,22,36,35,19,1,2,2,0,0,45,42,55,55,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,6,5,5,2,1,0,0,2,2,1,21,22,35,35,22,22,35,35,1,2,2,0,0,1,2,5,5,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,55,5,46,1,0,0,2,2,1,36,22,35,35,22,22,35,19,1,2,2,0,0,2,46,55,55,5,37,1,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,2,23,23,1,1,1,1,1,1,1,23,23,2,0,0,0,0,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,2,23,2,1,1,1,1,1,1,1,23,23,2,0,0,0,0,2,1,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,23,23,23,2,2,2,2,2,2,2,23,23,2,0,0,0,0,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,21,36,21,21,36,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,36,21,36,36,36,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,23,36,22,21,21,21,36,21,21,36,21,22,36,23,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,23,22,21,23,21,22,21,36,23,21,22,36,23,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,23,22,21,23,21,22,21,23,23,21,22,23,23,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,21,22,23,2,23,21,22,21,23,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,22,22,2,2,2,2,22,22,21,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,22,36,22,22,23,2,2,23,22,22,36,22,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,21,36,23,23,23,0,0,0,0,23,36,23,36,21,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,46,39,44,39,42,2,0,0,0,0,2,42,39,44,39,46,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,42,14,14,14,15,2,0,0,0,0,2,15,14,14,14,42,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,42,14,14,14,15,2,0,0,0,0,2,15,14,14,14,42,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,45,46,0,0,0,0,0,0,0,0,46,45,46,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0}
};



powerhero_text <=
'{
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,42,2,1,45,46,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,42,2,1,45,46,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,1,46,43,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,46,46,46,45,1,1,1,42,15,46,46,46,46,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,46,45,46,46,46,42,45,1,1,1,42,15,46,45,46,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,43,46,2,2,15,42,1,1,1,2,2,42,43,46,46,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,2,1,15,42,1,2,15,43,46,2,1,1,1,43,43,46,46,46,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,46,46,2,2,15,42,1,1,46,46,46,2,1,1,1,43,43,46,46,46,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,46,42,15,46,1,1,1,2,2,46,2,1,1,45,46,43,46,45,2,2,43,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,46,42,15,46,1,1,1,1,2,42,2,1,1,1,46,15,42,46,1,1,15,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,1,45,46,15,46,1,1,1,1,2,46,2,1,1,1,46,15,42,46,1,2,43,43,46,46,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,1,2,15,43,42,46,43,43,43,15,42,1,2,15,42,1,2,15,43,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,1,2,15,15,42,45,43,43,43,43,42,1,2,24,43,1,2,15,15,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,46,46,43,43,2,2,43,43,42,42,19,19,19,19,15,45,2,2,45,1,45,15,43,43,46,2,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,43,43,15,43,45,42,43,8,49,49,49,49,49,49,40,1,45,46,43,43,46,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,15,15,15,43,45,46,42,38,49,49,49,49,49,49,39,1,2,45,43,15,42,46,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,43,43,43,15,19,33,33,49,49,49,49,49,49,49,8,19,19,19,15,43,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,45,42,45,19,49,49,49,49,49,14,44,44,14,49,49,49,49,49,19,45,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,1,2,46,43,43,46,42,2,15,49,49,49,49,49,26,44,44,26,49,49,49,49,49,15,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,43,46,42,33,41,49,49,49,49,50,14,52,52,14,50,49,49,49,49,41,33,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,46,42,49,49,49,49,49,50,44,52,52,52,52,44,50,49,49,49,49,49,15,45,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,15,46,42,49,49,49,49,49,50,44,52,52,52,52,44,50,49,49,49,49,49,42,45,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,46,43,43,2,45,49,49,49,49,8,50,26,14,14,14,14,26,50,8,49,49,49,49,45,2,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,46,46,45,43,43,1,2,49,49,49,8,27,50,50,14,44,44,14,50,50,27,8,49,49,49,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,46,46,45,42,42,1,2,49,49,49,49,50,50,50,14,44,44,14,50,50,50,25,49,49,49,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,33,39,45,45,42,33,50,50,50,50,50,50,27,27,50,50,50,50,50,50,39,42,45,45,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,40,38,42,45,1,13,50,50,50,50,50,50,50,50,50,50,50,50,50,50,44,1,45,42,41,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,45,33,40,42,45,1,13,50,50,50,50,50,50,50,50,50,50,50,50,50,50,44,1,45,42,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,39,39,45,45,33,47,3,12,45,42,42,42,42,42,42,15,42,45,12,3,48,33,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,40,45,45,39,38,7,12,1,2,45,45,45,45,2,45,2,1,12,7,38,39,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,39,45,45,39,38,7,12,1,45,45,45,45,45,45,45,45,1,12,7,48,39,45,45,39,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,55,55,7,12,1,37,55,54,54,54,54,55,37,1,12,3,55,55,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,55,5,7,12,1,37,55,54,55,55,54,55,37,1,12,7,55,55,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,54,55,3,12,2,47,55,54,54,54,54,55,37,2,12,3,54,54,2,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,45,45,1,43,55,54,55,55,55,55,54,54,54,55,54,54,54,54,42,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,45,45,2,15,55,55,55,55,54,55,55,55,55,54,54,54,54,55,15,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,42,38,38,38,54,55,38,38,38,38,55,54,38,48,38,42,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,1,1,45,44,48,55,33,44,44,33,55,48,44,13,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,1,1,1,46,39,38,55,39,44,44,39,55,38,39,42,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,15,15,19,15,15,24,37,15,15,15,15,37,24,15,15,13,15,15,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,2,46,50,50,49,33,1,1,1,2,45,45,2,1,1,1,44,52,27,50,46,2,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,1,2,50,50,49,33,1,1,1,2,45,46,2,1,1,1,44,52,27,50,2,1,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,24,33,24,33,19,33,33,33,33,40,41,44,44,33,33,33,44,13,14,14,39,37,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,1,1,38,38,23,23,1,19,49,49,49,49,49,52,14,49,49,49,19,1,44,52,17,38,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,1,1,1,40,38,23,23,1,33,49,49,49,49,49,52,14,49,49,49,33,1,10,52,17,38,1,1,1,0,0,0,0,0,0},
'{0,0,0,0,0,24,54,33,15,47,48,2,2,0,0,42,8,49,50,14,8,49,49,8,42,0,0,13,13,38,38,33,33,54,24,0,0,0,0,0},
'{0,0,0,0,1,37,6,48,39,47,48,2,0,0,0,1,39,49,52,52,49,49,49,39,1,0,0,0,2,38,38,48,38,6,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,40,39,48,48,2,0,0,0,1,40,49,14,52,49,49,49,40,1,0,0,0,2,38,38,39,47,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,55,55,42,2,0,0,2,2,1,44,14,8,49,49,49,50,39,1,2,2,0,0,45,42,55,55,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,6,5,5,2,1,0,0,2,2,1,44,52,49,49,49,49,50,44,1,2,2,0,0,1,2,5,5,5,37,1,0,0,0,0},
'{0,0,0,0,1,37,5,55,5,46,1,0,0,2,2,1,44,52,8,49,49,49,50,44,1,2,2,0,0,2,46,55,55,5,37,1,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,2,23,23,1,2,2,2,2,1,1,23,23,2,0,0,0,0,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,2,23,23,1,1,1,1,1,1,1,23,23,2,0,0,0,0,2,1,1,0,0,0,0,0,0},
'{0,0,0,0,0,0,2,2,2,0,0,0,0,2,23,23,23,2,2,2,2,2,2,2,23,23,2,0,0,0,0,2,2,2,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,21,36,21,21,36,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,36,21,36,36,36,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,23,36,22,21,21,21,36,21,21,36,21,22,36,23,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,23,22,21,23,21,22,21,36,23,21,22,36,23,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,23,22,21,23,21,22,21,23,23,21,22,23,23,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,23,21,22,23,2,23,21,22,21,23,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,21,36,22,22,2,2,2,2,22,22,21,21,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,22,22,36,22,22,23,2,2,23,22,22,36,22,22,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,23,21,36,23,23,23,0,0,0,0,23,36,23,36,21,23,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,2,2,23,23,23,2,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,46,39,44,39,42,2,0,0,0,0,2,42,39,44,39,46,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,42,14,14,14,15,2,0,0,0,0,2,15,14,14,14,42,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,2,42,14,14,14,15,2,0,0,0,0,2,15,14,14,14,42,2,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,46,45,46,0,0,0,0,0,0,0,0,46,45,46,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0}
};

end

always_comb
begin
if (change ==1 )
hero_text=powerhero_text;

else
hero_text=hero123_text	;
end


endmodule
